`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Long Chen
// Create Date: 2023/11/30 19:18:12
// Design Name: enigma_top
// Module Name:  enigma_top
// Project Name: ENIGMA551
//////////////////////////////////////////////////////////////////////////////////


module enigma_top(

    );
endmodule
