`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/30/2023 11:45:54 PM
// Design Name: 
// Module Name: enigma_onward_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module enigma_onward_sim(

    );
    
reg rst;
reg [4:0]data_in;
wire [4:0]data_out;
wire [4:0]r1;
wire [4:0]r2;
wire [4:0]r3;
wire [4:0]r11;
wire [4:0]r22;
wire [4:0]r33;
integer i;
initial
begin
rst=1'd0;
data_in=5'd0;
end
enigma_implementation_onward eio(.rst(rst),.data_in(data_in),.data_out(data_out),
.r1_positionF(r1),.r2_positionF(r2),.r3_positionF(r3),
.r1_positionB(r11),.r2_positionB(r22),.r3_positionB(r33));
initial
begin

for(i=0;i<5000;i=i+1)begin
if(data_in==5'd25)begin
data_in=5'd0;
end
else
begin
 data_in=data_in+5'd1;
 end
 #5;
 end
/*
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
*/
/*
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
#1 data_in=5'd0;
#1 data_in=5'd1;
#1 data_in=5'd2;
#1 data_in=5'd3;
#1 data_in=5'd4;
#1 data_in=5'd5;
#1 data_in=5'd6;
#1 data_in=5'd7;
#1 data_in=5'd8;
#1 data_in=5'd9;
#1 data_in=5'd10;
#1 data_in=5'd11;
#1 data_in=5'd12;
#1 data_in=5'd13;
#1 data_in=5'd14;
#1 data_in=5'd15;
#1 data_in=5'd16;
#1 data_in=5'd17;
#1 data_in=5'd18;
#1 data_in=5'd19;
#1 data_in=5'd20;
#1 data_in=5'd21;
#1 data_in=5'd22;
#1 data_in=5'd23;
#1 data_in=5'd24;
#1 data_in=5'd25;
*/
end
endmodule
